** Copyright: Suming Lai
** Oct. 10, 2011
** Modified by: Honghuang Lin
** Sep. 10, 2015

.PARAM voutac=0 vdddc=1.2 vddac=0 il=0.000000e+00 ib=5u cf=1.600000e-13 cz=2.000000e-13 cc2=4.000000e-13 cc1=1.000000e-12 Rf1=7.800000e+04 Rf2=1.220000e+05

**.AC DEC 200 1.000000e+00 1.000000e+12

.TRAN 1n 16u

.TEMP 25
.OPTION
+    ARTIST=2
+    INGOLD=2
+    MEASOUT=1
+    PARHIER=LOCAL
+    POST
+    PSF=2
+    NOMOD
+        MEASDGT=7
* set the measure output digits

.inc ./param0.inc
.INCLUDE "../tech/hspice.include"
.inc ../tech/nfet_perfect.inc
.inc ../tech/pfet_perfect.inc

ib vbias2x my_gnd DC=ib

cz vfb2x vout cz
c2 ampoutpx my_gnd cc2
c1 amp1outpx my_gnd cc1
cc ampoutpx vfb2x cf
r1 vout vfb2x Rf1
r2 vfb2x my_gnd Rf2
iLoad vout 0 PWL 0 0.005 1u 0.005 1.1u 0.105 3u 0.105

v0 my_gnd 0 DC=0 AC=0

vr vref2 0 DC=610e-3 AC=0

vcc my_vdd 0 DC=vdddc AC=vddac

** M1
xt1 net0237 ampoutpx vout vout pfet l='80e-9+l7*920e-9' w='120e-9+w7*49880e-9' par=1 m=1 nf=200 dtemp=0 rgatemod=0 sa=240e-9 sb=240e-9 sd=280e-9 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 lmlt=1 vmlt=1 omlt=1

** M2
xt2 net0237 amp1outnx my_gnd my_gnd nfet l='8.000000e-08' w=2.700000e-05 par=1 m=1 nf=30 ptwell=1 dtemp=0 rgatemod=0 sa=240e-9 sb=240e-9 sd=280e-9 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 lmlt=1 vmlt=1 omlt=1

** M3
xt3 amp1outpx vref2 net0167 net0167 pfet l='80e-9+l1*920e-9' w='120e-9+w1*49880e-9' par=1 ad=1.92e-12 as=2.12e-12 pd=15.84e-6 ps=18.24e-6 m=1 nf=12 dtemp=0 rgatemod=0 sa=260e-9 sb=260e-9 sd=320e-9 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 lmlt=1 vmlt=1 omlt=1

** M4
xt4 amp1outnx vfb2x net0167 net0167 pfet l='80e-9+l2*920e-9' w='120e-9+w2*49880e-9' par=1 ad=1.92e-12 as=2.12e-12 pd=15.84e-6 ps=18.24e-6 m=1 nf=12 dtemp=0 rgatemod=0 sa=260e-9 sb=260e-9 sd=320e-9 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 lmlt=1 vmlt=1 omlt=1

** M6
xt5 amp1outpx vref2 net0278 my_gnd nfet l='80e-9+l3*920e-9' w='120e-9+w3*49880e-9' par=1 ad=153.6e-15 as=201.6e-15 pd=2.24e-6 ps=3.12e-6 m=1 nf=4 ptwell=1 dtemp=0 rgatemod=0 sa=260e-9 sb=260e-9 sd=320e-9 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 lmlt=1 vmlt=1 omlt=1

** M5
xt6 amp1outnx vfb2x net0278 my_gnd nfet l='80e-9+l4*920e-9' w='120e-9+w4*49880e-9' par=1 ad=153.6e-15 as=201.6e-15 pd=2.24e-6 ps=3.12e-6 m=1 nf=4 ptwell=1 dtemp=0 rgatemod=0 sa=260e-9 sb=260e-9 sd=320e-9 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 lmlt=1 vmlt=1 omlt=1

** M7
xt7 amp1outpx amp1outpx my_gnd my_gnd nfet l='160e-9' w=700e-9 par=1 ad=112e-15 as=147e-15 pd=1.98e-6 ps=2.73e-6 m=1 nf=4 ptwell=1 dtemp=0 rgatemod=0 sa=260e-9 sb=260e-9 sd=320e-9 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 lmlt=1 vmlt=1 omlt=1

** M8
xt8 amp1outnx amp1outnx my_gnd my_gnd nfet l='160e-9' w=700e-9 par=1 ad=112e-15 as=147e-15 pd=1.98e-6 ps=2.73e-6 m=1 nf=4 ptwell=1 dtemp=0 rgatemod=0 sa=260e-9 sb=260e-9 sd=320e-9 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 lmlt=1 vmlt=1 omlt=1

** M9
xt9 amp1outpx amp1outnx my_gnd my_gnd nfet l='80e-9+l5*920e-9' w='120e-9+w5*49880e-9' par=1 ad=105.6e-15 as=138.6e-15 pd=1.94e-6 ps=2.67e-6 m=1 nf=4 ptwell=1 dtemp=0 rgatemod=0 sa=260e-9 sb=260e-9 sd=320e-9 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 lmlt=1 vmlt=1 omlt=1

** M10
xt10 amp1outnx amp1outpx my_gnd my_gnd nfet l='80e-9+l6*920e-9' w='120e-9+w6*49880e-9' par=1 ad=105.6e-15 as=138.6e-15 pd=1.94e-6 ps=2.67e-6 m=1 nf=4 ptwell=1 dtemp=0 rgatemod=0 sa=260e-9 sb=260e-9 sd=320e-9 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 lmlt=1 vmlt=1 omlt=1

** M11
xt11 ampoutpx amp1outpx my_gnd my_gnd nfet l='120e-9' w=2.2e-6 par=1 ad=352e-15 as=572e-15 pd=2.84e-6 ps=5.44e-6 m=1 nf=2 ptwell=1 dtemp=0 rgatemod=0 sa=260e-9 sb=260e-9 sd=320e-9 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 lmlt=1 vmlt=1 omlt=1

** M12
xtp1 vout net0237 my_vdd my_vdd pfet l='80e-9' w=4.500000e-04 par=1 m=1 nf=500 dtemp=0 rgatemod=0 sa=240e-9 sb=240e-9 sd=280e-9 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 lmlt=1 vmlt=1 omlt=1

** M13
xtpn vout net0237 my_gnd my_gnd nfet l='80e-9+l8*920e-9' w='120e-9+w8*49880e-9' par=1 ad=117e-15 as=117e-15 pd=1.42e-6 ps=1.42e-6 m=1 nf=1 ptwell=1 dtemp=0 rgatemod=0 sa=260e-9 sb=260e-9 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 lmlt=1 vmlt=1 omlt=1

** M14
xtb0 vbias2x vbias2x my_vdd my_vdd pfet l='960e-9' w=9.6e-6 par=1 ad=1.536e-12 as=2.016e-12 pd=10.88e-6 ps=16.08e-6 m=1 nf=4 dtemp=0 rgatemod=0 sa=260e-9 sb=260e-9 sd=320e-9 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 lmlt=1 vmlt=1 omlt=1

** M15
xtb1 net0183 vbias2x my_vdd my_vdd pfet l='960e-9' w=9.6e-6 par=1 ad=1.536e-12 as=2.016e-12 pd=10.88e-6 ps=16.08e-6 m=1 nf=4 dtemp=0 rgatemod=0 sa=260e-9 sb=260e-9 sd=320e-9 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 lmlt=1 vmlt=1 omlt=1

** M16
xtb2 net0167 vbias2x my_vdd my_vdd pfet l='960e-9' w=96e-6 par=1 ad=15.36e-12 as=15.84e-12 pd=108.8e-6 ps=114e-6 m=1 nf=40 dtemp=0 rgatemod=0 sa=260e-9 sb=260e-9 sd=320e-9 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 lmlt=1 vmlt=1 omlt=1

** M17
xtb3 ampoutpx vbias2x my_vdd my_vdd pfet l='960e-9' w=14.4e-6 par=1 ad=2.304e-12 as=2.784e-12 pd=16.32e-6 ps=21.52e-6 m=1 nf=6 dtemp=0 rgatemod=0 sa=260e-9 sb=260e-9 sd=320e-9 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 lmlt=1 vmlt=1 omlt=1

** M18
xtbn0 net0278 vbias1x my_gnd my_gnd nfet l='480e-9' w=6e-6 par=1 ad=960e-15 as=1.02e-12 pd=12.4e-6 ps=13.4e-6 m=1 nf=20 ptwell=1 dtemp=0 rgatemod=0 sa=260e-9 sb=260e-9 sd=320e-9 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 lmlt=1 vmlt=1 omlt=1

** M19
xtbn1 vbias1x vbias1x my_gnd my_gnd nfet l='480e-9' w=1.2e-6 par=1 ad=192e-15 as=252e-15 pd=2.48e-6 ps=3.48e-6 m=1 nf=4 ptwell=1 dtemp=0 rgatemod=0 sa=260e-9 sb=260e-9 sd=320e-9 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 lmlt=1 vmlt=1 omlt=1

** M20
xtbn2 vbias1x vbias1x net0183 net0183 pfet l='480e-9' w=9.6e-6 par=1 ad=1.536e-12 as=2.016e-12 pd=10.88e-6 ps=16.08e-6 m=1 nf=4 dtemp=0 rgatemod=0 sa=260e-9 sb=260e-9 sd=320e-9 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=0 panw10=0 lmlt=1 vmlt=1 omlt=1

*.ALTER
*.param0  voutac=1 vddac=0
.OP

.MEAS TRAN iq0 AVG I(vcc) FROM=0u TO=0.1u
.MEAS TRAN iq1 AVG I(vcc) FROM=15.9u TO=16u
.MEAS TRAN uds MIN V(vout) FROM=0u TO=6u
.MEAS TRAN vout0 AVG V(vout) FROM=0n TO=100n
.MEAS TRAN vout1 AVG V(vout) FROM=15.9u TO=16u
.MEAS TRAN voutr AVG V(vout) FROM=15.8u TO=15.9u